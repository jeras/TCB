////////////////////////////////////////////////////////////////////////////////
// TCB peripheral: UART controller package
////////////////////////////////////////////////////////////////////////////////
// Copyright 2022 Iztok Jeras
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
////////////////////////////////////////////////////////////////////////////////

module tcb_peri_uart_pkg;

    // helper function for calculating boudrate divider
    function int unsigned baudrate_divider (
        input  int unsigned frequency,          // Hz units
        input  int unsigned baudrate = 115200   // Hz units
    );
        return frequency/baudrate;
    endfunction: baudrate_divider

endmodule: tcb_peri_uart_pkg
