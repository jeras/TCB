////////////////////////////////////////////////////////////////////////////////
// TCB interface UART controller, asynchronous deserializer
////////////////////////////////////////////////////////////////////////////////
// Copyright 2022 Iztok Jeras
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
////////////////////////////////////////////////////////////////////////////////

module tcb_uart_des #(
  int unsigned CW = 8,  // baudrate counter width
  int unsigned DW = 8   // shifter data width
)(
  // system signals
  input  logic          clk,
  input  logic          rst,
  // configuration
  input  logic [CW-1:0] cfg_bdr,  // baudrate
  input  logic [CW-1:0] cfg_smp,  // sample position
  // parallel stream (there is no READY signal)
  output logic          str_vld,  // valid
  output logic [DW-1:0] str_dat,  // data
  // serial RX output
  input  logic          rxd
);

// parallel stream transfer
logic          str_trn;

// baudrate counter
logic [CW-1:0] bdr_cnt;
logic          bdr_end;
logic          bdr_hlf;

// shifter bit counter
logic  [4-1:0] shf_cnt;
logic  [4-1:0] shf_end;

// shift data register
logic [DW-1:0] shf_dat;

// delay RDX and detect a start edge
logic          rxd_dly;
logic          rxd_edg;

////////////////////////////////////////////////////////////////////////////////
// parallel stream
////////////////////////////////////////////////////////////////////////////////

// parallel stream transfer
assign str_trn = str_vld;

// parallel stream valid
assign str_vld = shf_end;

////////////////////////////////////////////////////////////////////////////////
// start bit detection
////////////////////////////////////////////////////////////////////////////////

// delay uart_rxd and detect a start negative edge
always @ (posedge clk)
rxd_dly <= rxd;

assign rxd_start = rxd_dly & ~rxd;

////////////////////////////////////////////////////////////////////////////////
// serializer
////////////////////////////////////////////////////////////////////////////////

// baudrate generator from clock (it counts down to 0 generating a baud pulse)
always @ (posedge clk, posedge rst)
if (rst)        bdr_cnt <= '0;
else begin
  if (str_trn)  bdr_cnt <= '0;
  else          bdr_cnt <= bdr_cnt + (~shf_end);
end

// enable signal for shifting logic
assign bdr_end = bdr_cnt == cfg_bdr;

// enable signal for sample logic
assign bdr_smp = bdr_cnt == cfg_smp;

// bit counter
always @ (posedge clk, posedge rst)
if (rst)        shf_cnt <= 4'd0;
else begin
  if (str_trn)  shf_cnt <= 4'(DW);
  else          shf_cnt <= shf_cnt - 1;
end

// end of shift sequence
assign shf_end = shf_cnt == 4'd0;

// data shift register
always @ (posedge clk)
if (bdr_smp)  shf_dat <= {rxd, shf_dat[DW-1:1]};

// parallel stream data
assign str_dat = shf_dat;

endmodule: tcb_uart_des