////////////////////////////////////////////////////////////////////////////////
// TCB-Lite peripheral: GPIO controller
//
// NOTE: In case this module is connected to asynchronous signals,
//       the input signals `gpio_i` require a CDC synchronizer.
//       By default a 2 FF synchronizer is implemented by the CFG_CDC parameter.
////////////////////////////////////////////////////////////////////////////////
// Copyright 2023 Iztok Jeras
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
////////////////////////////////////////////////////////////////////////////////

module tcb_lite_peri_gpio #(
    // GPIO parameters
    parameter  int unsigned GDW = 32,  // GPIO data width
    parameter  int unsigned CDC =  2,  // implement clock domain crossing stages (0 - bypass)
    // optional implementation configuration
    parameter  bit           CFG_IEN =   '0,  // input enable implementation
    parameter  bit [GDW-1:0] CFG_IRQ =   '1,  // interrupt request implementation mask
    parameter  bit           CFG_MIN = 1'b0   // minimalistic response implementation (configuration is write only)
    // NOTE 1: if none of the interrupts are enabled, the controller has a smaller address space
)(
    // GPIO signals
    output logic [GDW-1:0] gpio_o,
    output logic [GDW-1:0] gpio_e,
    input  logic [GDW-1:0] gpio_i,
    // TCB interface
    tcb_lite_if.sub sub,
    // IRQ interface
    output logic irq
);

////////////////////////////////////////////////////////////////////////////////
// parameter validation
////////////////////////////////////////////////////////////////////////////////

    initial begin
        assert (sub.DLY ==   0) else $error("unsupported DLY = %0d (must be 0)", sub.DLY);
        assert (sub.DAT >= GDW) else $error("unsupported (DAT = %0d) < (GDW = %0d)", sub.DAT, GDW);
    end

////////////////////////////////////////////////////////////////////////////////
// GPIO instance
////////////////////////////////////////////////////////////////////////////////

    logic [3-1:0] sys_req_adr;

    // check whether at least one GPIO pin has enabled interrupt support
    generate
    if (~CFG_IRQ) begin
        assign sys_req_adr =        sub.req.adr[sub.MAX+:3];
    end else begin
        assign sys_req_adr = {1'b0, sub.req.adr[sub.MAX+:2]};
    end
    endgenerate


    tcb_peri_gpio #(
        // GPIO parameters
        .GDW      (GDW),
        .CDC      (CDC),
        // system interface parameters
        .DAT      (sub.DAT),
        // optional implementation configuration
        .CFG_IEN  (CFG_IEN),
        .CFG_IRQ  (CFG_IRQ),
        .CFG_MIN  (CFG_MIN)
    ) gpio (
        // GPIO signals
        .gpio_o   (gpio_o),
        .gpio_e   (gpio_e),
        .gpio_i   (gpio_i),
        // system signals
        .clk      (sub.clk),
        .rst      (sub.rst),
        // system write interface
        .sys_wen  (sub.req.wen & sub.trn),
        .sys_wad  (sys_req_adr),
        .sys_wdt  (sub.req.wdt),
        // system read interface
        .sys_ren  (~sub.req.wen & sub.trn),
        .sys_rad  (sys_req_adr),
        .sys_rdt  (sub.rsp.rdt),
        // interrupt request interface
        .irq      (irq)
    );

    // status response
    assign sub.rsp.sts =   '0;
    assign sub.rsp.err = 1'b0;

endmodule: tcb_lite_peri_gpio
