////////////////////////////////////////////////////////////////////////////////
// SPI slave model
////////////////////////////////////////////////////////////////////////////////
// Copyright 2025 Iztok Jeras
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
////////////////////////////////////////////////////////////////////////////////

module spi_slave_model
    import spi_pkg::*;
#(
    // shift register width
    parameter  int unsigned DAT = 8,
    // IO data width (supported values are 2, 4, 8)
    parameter  int unsigned IO_WIDTH = 2
)(
    input  wire                sclk,  // serial clock
    input  wire                ss_n,  // slave select
    inout  wire [IO_WIDTH-1:0] sdio   // serial data I/O {sdio[IO_WIDTH-1:2], miso, mosi}
);

endmodule: spi_slave_model
