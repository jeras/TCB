////////////////////////////////////////////////////////////////////////////////
// TCB-Lite (Tightly Coupled Bus) library demultiplexer/decoder testbench
////////////////////////////////////////////////////////////////////////////////
// Copyright 2022 Iztok Jeras
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
////////////////////////////////////////////////////////////////////////////////

module tcb_lite_lib_demultiplexer_tb
    import tcb_lite_pkg::*;
#(
    // RTL configuration parameters
    parameter  int unsigned DLY =    1,  // response delay
    parameter  bit          HLD = 1'b0,  // response hold
    parameter  bit          MOD = 1'b1,  // bus mode (0-logarithmic size, 1-byte enable)
    parameter  int unsigned CTL =    0,  // control width (user defined request signals)
    parameter  int unsigned ADR =   32,  // address width (only 32/64 are supported)
    parameter  int unsigned DAT =   32,  // data    width (only 32/64 are supported)
    parameter  int unsigned STS =    0,  // status  width (user defined response signals)
    // interconnect parameters (interface number)
    parameter  int unsigned IFN = 3,
    localparam int unsigned IFL = $clog2(IFN)
);

////////////////////////////////////////////////////////////////////////////////
// local parameters
////////////////////////////////////////////////////////////////////////////////

    // decoder address and mask array
    localparam logic [ADR-1:0] DAM [IFN-1:0] = '{
        ADR'({14'bx, 2'b1x, 16'hxxxx}),
        ADR'({14'bx, 2'b01, 16'hxxxx}),
        ADR'({14'bx, 2'b00, 16'hxxxx})
    };

    // TCB configurations               '{HSK: '{DLY, HLD}, BUS: '{MOD, CTL, ADR, DAT, STS}}
    localparam tcb_lite_cfg_t MAN_CFG = '{HSK: '{DLY, HLD}, BUS: '{MOD, CTL, ADR, DAT, STS}};
    localparam tcb_lite_cfg_t SUB_CFG = '{HSK: '{DLY, HLD}, BUS: '{MOD, CTL, ADR, DAT, STS}};

    localparam bit VIP = 1'b1;

////////////////////////////////////////////////////////////////////////////////
// local signals
////////////////////////////////////////////////////////////////////////////////

    // system signals (initialized)
    logic clk = 1'b1;  // clock
    logic rst = 1'b1;  // reset

    string testname = "none";

    // TCB interfaces
    tcb_lite_if #(MAN_CFG) tcb_man           (.clk (clk), .rst (rst));
    tcb_lite_if #(SUB_CFG) tcb_sub [IFN-1:0] (.clk (clk), .rst (rst));

    // empty array
    logic [8-1:0] nul [];

    // response
    logic [DAT-1:0] rdt;  // read data
    logic [STS-1:0] sts;  // response status
    logic           err;  // response error

    // control
    logic [IFL-1:0] sel;  // select

////////////////////////////////////////////////////////////////////////////////
// tests
////////////////////////////////////////////////////////////////////////////////

    task test_simple ();
        // write sequence
        $display("write sequence");
//        testname = "write";
//        for (int i=0; i<IFN; i++) begin
//            tst_sub[i].delete();
//            tst_mon[i].delete();
//        end
//        fork
//            // manager (blocking API)
//            begin: fork_man
//                for (int unsigned i=0; i<IFN; i++) begin
//                    obj_man.write32((i<<16) + 32'h00000000, 32'h76543210, sts);
//                    obj_man.write32((i<<16) + 32'h00000020, 32'hfedcba98, sts);
//                    obj_man.read32 ((i<<16) + 32'h00000000, rdt[4-1:0], sts);
//                    obj_man.read32 ((i<<16) + 32'h00000020, rdt[4-1:0], sts);
//                end
//            end: fork_man
//            // subordinate (driver)
//            for (int unsigned i=0; i<IFN; i++)
//            begin: fork_sub_driver
//                sts[i] = '0;
//                tst_len[i] = tst_sub[i].size();
//                // append reference transfers to queue                        adr                wdt
//                tst_len[i] += obj_sub[i].put_transaction(tst_sub[i], '{req: '{adr: 32'h00000000, wdt: '{8'h10, 8'h32, 8'h54, 8'h76}, default: 'x}, rsp: '{nul, sts}});
//                tst_len[i] += obj_sub[i].put_transaction(tst_sub[i], '{req: '{adr: 32'h00000020, wdt: '{8'h98, 8'hba, 8'hdc, 8'hfe}, default: 'x}, rsp: '{nul, sts}});
//                tst_len[i] += obj_sub[i].put_transaction(tst_sub[i], '{req: '{adr: 32'h00000000, wdt: nul, default: 'x}, rsp: '{'{8'h10, 8'h32, 8'h54, 8'h76}, sts}});
//                tst_len[i] += obj_sub[i].put_transaction(tst_sub[i], '{req: '{adr: 32'h00000020, wdt: nul, default: 'x}, rsp: '{'{8'h98, 8'hba, 8'hdc, 8'hfe}, sts}});
////                for (int unsigned j=0; j<tst_sub[i].size(); j++) begin
////                  $display("DEBUG: tst_sub[%0d][%0d] = %p", i, j, tst_sub[i][j]);
////                end
//                obj_sub[i].transfer_sequencer(tst_sub[i]);
//            end: fork_sub_driver
//            // subordinate (monitor)
//            for (int unsigned i=0; i<IFN; i++)
//            begin: fork_sub_monitor
//                obj_sub[i].transfer_monitor(tst_mon[i]);
//            end: fork_sub_monitor
//        join_any
//        // disable transfer monitor
//        repeat (tcb_man.CFG.HSK.DLY) @(posedge clk);
//        disable fork;
//        // reference transfer queue
//        for (int unsigned i=0; i<IFN; i++)
//        begin
//            // compare transfers from monitor to reference
//            // wildcard operator is used to ignore data byte comparison, when the reference data is 8'hxx
//            for (int unsigned j=0; j<tst_sub[i].size(); j++) begin
//                assert (tst_mon[i][j].req ==? tst_sub[i][j].req) else $error("\ntst_mon[%0d][%0d].req = %p !=? \ntst_sub[%0d][%0d].req = %p", i, j, tst_mon[i][j].req, i, j, tst_sub[i][j].req);
//                assert (tst_mon[i][j].rsp ==? tst_sub[i][j].rsp) else $error("\ntst_mon[%0d][%0d].rsp = %p !=? \ntst_sub[%0d][%0d].rsp = %p", i, j, tst_mon[i][j].rsp, i, j, tst_sub[i][j].rsp);
//            end
////            // printout transfer queue for debugging purposes
////            for (int unsigned j=0; j<tst_sub[i].size(); j++) begin
////              $display("DEBUG: tst_sub[%0d][%0d] = %p", i, j, tst_sub[i][j]);
////              $display("DEBUG: tst_mon[%0d][%0d] = %p", i, j, tst_mon[i][j]);
////            end
//        end
    endtask: test_simple

////////////////////////////////////////////////////////////////////////////////
// test sequence
////////////////////////////////////////////////////////////////////////////////

    // clock
    always #(20ns/2) clk = ~clk;

    // test sequence
    initial
    begin: test
        // reset sequence
        repeat (2) @(posedge clk);
        /* verilator lint_off INITIALDLY */
        rst <= 1'b0;
        /* verilator lint_on INITIALDLY */
        repeat (1) @(posedge clk);

        test_simple;
//        test_parameterized;

        // end of test
        repeat (4) @(posedge clk);
        $finish();
    end: test

////////////////////////////////////////////////////////////////////////////////
// VIP instances
////////////////////////////////////////////////////////////////////////////////

    // manager VIP
    tcb_lite_vip_manager #(
    ) man (
        .man (tcb_man)
    );

    // subordinate VIP
    tcb_lite_vip_subordinate #(
    ) sub [IFN-1:0] (
        .sub (tcb_sub)
    );

    // manager TCB-Lite protocol checker
    tcb_lite_vip_protocol_checker chk_man (
        .mon (tcb_man)
    );

    // subordinate TCB-Lite protocol checker
    tcb_lite_vip_protocol_checker chk_sub [IFN-1:0] (
        .mon (tcb_sub)
    );

////////////////////////////////////////////////////////////////////////////////
// DUT instances
////////////////////////////////////////////////////////////////////////////////

    // RTL decoder DUT
    tcb_lite_lib_decoder #(
        // interconnect parameters
        .IFN  (IFN),
        // decoder address and mask array
        .DAM  (DAM)
    ) dut_dec (
        .mon  (tcb_man),
        .sel  (sel)
    );

    // RTL demultiplexer DUT
    tcb_lite_lib_demultiplexer #(
        // interconnect parameters
        .IFN   (IFN)
    ) dut_dmx (
        // control
        .sel  (sel),
        // TCB interfaces
        .sub  (tcb_man),
        .man  (tcb_sub)
    );

////////////////////////////////////////////////////////////////////////////////
// VCD/FST waveform trace
////////////////////////////////////////////////////////////////////////////////

    initial
    begin
`ifdef VERILATOR
        $dumpfile("test.fst");
`else
        $dumpfile("test.vcd");
`endif
        $dumpvars;
    end

endmodule: tcb_lite_lib_demultiplexer_tb
