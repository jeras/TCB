////////////////////////////////////////////////////////////////////////////////
// SPI master model
////////////////////////////////////////////////////////////////////////////////
// Copyright 2025 Iztok Jeras
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
////////////////////////////////////////////////////////////////////////////////

module spi_master_model
    import spi_pkg::*;
#(
    // default clock period
    parameter  realtime     PERIOD = 20ns,  // 50MHz
    // IO data width (supported values are 2, 4, 8)
    parameter  int unsigned IO_WIDTH = 2
)(
    inout  wire                sclk,  // serial clock
    output wire                ss_n,  // slave select
    inout  wire [IO_WIDTH-1:0] sdio   // serial data I/O {sdio[IO_WIDTH-1:2], miso, mosi}
);

////////////////////////////////////////////////////////////////////////////////
// local configuration accessible from outside
////////////////////////////////////////////////////////////////////////////////

    // clock period (initialized with parameter)
    realtime cfg_period = PERIOD;

    // SPI mode
    spi_mode_t cfg_mode = SPI_MODE0;

    // SPI width (single, dual, quad, octa)
    spi_width_e cfg_width = SPI_SINGLE;

    // SPI duplex (half, dual)
    spi_duplex_e cfg_duplex = SPI_FULL;

////////////////////////////////////////////////////////////////////////////////
// local signals
////////////////////////////////////////////////////////////////////////////////

    logic                clk;  // clock
    logic                sel;  // select
    logic                oen;  // output enable
    logic [IO_WIDTH-1:0] dti;  // data input
    logic [IO_WIDTH-1:0] dto;  // data output

////////////////////////////////////////////////////////////////////////////////
// initialization
////////////////////////////////////////////////////////////////////////////////


////////////////////////////////////////////////////////////////////////////////
// transaction
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// I/O
////////////////////////////////////////////////////////////////////////////////



endmodule: spi_master_model