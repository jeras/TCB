////////////////////////////////////////////////////////////////////////////////
// TCB-Lite (Tightly Coupled Bus) library register slice for request path
////////////////////////////////////////////////////////////////////////////////
// Copyright 2022 Iztok Jeras
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
////////////////////////////////////////////////////////////////////////////////

module tcb_lite_lib_register_request
    import tcb_lite_pkg::*;
#(
    parameter string OPT = "POWER"  // optimization for "POWER" or "COMPLEXITY"
)(
    // TCB-Lite interfaces
    tcb_lite_if.sub sub,  // TCB subordinate interface (manager     device connects here)
    tcb_lite_if.man man   // TCB manager     interface (subordinate device connects here)
);

////////////////////////////////////////////////////////////////////////////////
// parameter validation
////////////////////////////////////////////////////////////////////////////////

`ifdef ALTERA_RESERVED_QIS
`else
    // comparing subordinate and manager interface parameters
    initial
    begin
        assert (man.CFG.HSK.DLY+1 == sub.CFG.HSK.DLY) else $error("Parameter (man.CFG.HSK.DLY = %p)+1 != (sub.CFG.HSK.DLY = %p)", man.CFG.HSK.DLY, sub.CFG.HSK.DLY);

        assert (man.CFG.BUS == sub.CFG.BUS) else $error("Parameter (man.CFG.BUS = %p) != (sub.CFG.BUS = %p)", man.CFG.BUS, sub.CFG.BUS);
    end
`endif

////////////////////////////////////////////////////////////////////////////////
// register request path
////////////////////////////////////////////////////////////////////////////////

    // handshake
    always_ff @(posedge sub.clk, posedge sub.rst)
    if (sub.rst) begin
        man.vld <= 1'b0;
    end else begin
        if (sub.rdy) begin
            man.vld <= sub.vld;
        end
    end

    // request
    always_ff @(posedge sub.clk)
    if (sub.trn) begin
        man.req.lck <= sub.req.lck;
        man.req.wen <= sub.req.wen;
        man.req.ren <= sub.req.ren;
        man.req.ndn <= sub.req.ndn;
        man.req.ctl <= sub.req.ctl;
        man.req.adr <= sub.req.adr;
        man.req.siz <= sub.req.siz;
        man.req.byt <= sub.req.byt;
//        man.req.wdt <= sub.req.wdt;
    end

    generate
    case (OPT)
        "POWER": begin
            case (sub.CFG.BUS.MOD)
                // logarithmic size
                1'b0: begin: byt
                    // write data
                    for (genvar i=0; i<sub.CFG_BUS_BYT; i++) begin: wdt
                        always_ff @(posedge sub.clk)
                        if (sub.trn & sub.req.wen) begin
                            if (i < (1<<sub.req.siz)) begin
                                man.req.wdt[i*8+:8] <= sub.req.wdt[i*8+:8];
                            end
                        end
                    end: wdt
                end: byt
                // byte enable
                1'b1: begin: byt
                    // write data
                    for (genvar i=0; i<sub.CFG_BUS_BYT; i++) begin: wdt
                        always_ff @(posedge sub.clk)
                        if (sub.trn & sub.req.wen) begin
                            if (sub.req.byt[i]) begin
                                man.req.wdt[i*8+:8] <= sub.req.wdt[i*8+:8];
                            end 
                        end
                    end: wdt
                end: byt
            endcase
        end
        "COMPLEXITY": begin
            always_ff @(posedge sub.clk)
            if (sub.trn & sub.req.wen) begin
                man.req.wdt <= sub.req.wdt;
            end
        end
    endcase
    endgenerate

    // response
    assign sub.rsp.rdt = man.rsp.rdt;
    assign sub.rsp.sts = man.rsp.sts;
    assign sub.rsp.err = man.rsp.err;

    // handshake (valid is checked to avoid pipeline bubbles)
    assign sub.rdy = man.rdy | ~man.vld;

endmodule: tcb_lite_lib_register_request
